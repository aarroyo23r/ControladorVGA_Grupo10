`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/23/2017 03:14:40 PM
// Design Name: 
// Module Name: SelectorDeco
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module SelectorDeco(
    input [9:0] pixelx,
    input [9:0] pixely,
    output [6:0] Dir,
    input [6:0] Dir0,
    input [6:0] Dir1,
    input [6:0] Dir2,
    input [6:0] Dir3,
    input clock
    );
endmodule

// Bloque grande generador de datos
